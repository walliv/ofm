// property.sv
// Copyright (C) 2022-2024 CESNET z. s. p. o.
// Author(s): Daniel Kriz <danielkriz@cesnet.cz>
//            Vladislav Valek <valekv@cesnet.cz>

// SPDX-License-Identifier: BSD-3-Clause

import uvm_pkg::*;
`include "uvm_macros.svh"

module TX_DMA_CALYPTE_PROPERTY #(
    USR_TX_MFB_REGIONS,
    USR_TX_MFB_REGION_SIZE,
    USR_TX_MFB_BLOCK_SIZE,
    USR_TX_MFB_ITEM_WIDTH,

    USR_MFB_META_WIDTH,

    PCIE_CQ_MFB_REGIONS,
    PCIE_CQ_MFB_REGION_SIZE,
    PCIE_CQ_MFB_BLOCK_SIZE,
    PCIE_CQ_MFB_ITEM_WIDTH
) (
    input logic RESET,
    mfb_if cq_mfb,
    mfb_if usr_tx_mfb
);

    string module_name = "";
    logic START = 1'b1;

    ///////////////////
    // Start check properties after first clock
    initial begin
        $sformat(module_name, "%m");
        @(posedge usr_tx_mfb.CLK)
        #(10ps)
        START = 1'b0;
    end

    mfb_property #(
        .REGIONS     (PCIE_CQ_MFB_REGIONS                  ),
        .REGION_SIZE (PCIE_CQ_MFB_REGION_SIZE              ),
        .BLOCK_SIZE  (PCIE_CQ_MFB_BLOCK_SIZE               ),
        .ITEM_WIDTH  (PCIE_CQ_MFB_ITEM_WIDTH               ),
        .META_WIDTH  (sv_pcie_meta_pack::PCIE_CQ_META_WIDTH)
    ) cq_mfb_property_i (
        .RESET (RESET),
        .vif   (cq_mfb)
    );

    mfb_property #(
        .REGIONS     (USR_TX_MFB_REGIONS    ),
        .REGION_SIZE (USR_TX_MFB_REGION_SIZE),
        .BLOCK_SIZE  (USR_TX_MFB_BLOCK_SIZE ),
        .ITEM_WIDTH  (USR_TX_MFB_ITEM_WIDTH ),
        .META_WIDTH  (USR_MFB_META_WIDTH    )
    ) usr_tx_mfb_property_i (
        .RESET (RESET),
        .vif   (usr_tx_mfb)
    );
endmodule
